magic
tech sky130A
magscale 1 2
timestamp 1729052455
<< error_s >>
rect 54 2010 178 2023
rect 2031 2010 2125 2024
<< locali >>
rect -14 2556 2001 2575
rect -14 2508 83 2556
rect 1885 2508 2001 2556
rect -14 2492 2001 2508
rect 5 1501 2020 1518
rect 5 1453 32 1501
rect 1834 1453 2020 1501
rect 5 1435 2020 1453
<< viali >>
rect 83 2508 1885 2556
rect 32 1453 1834 1501
<< metal1 >>
rect -16 2556 2012 2575
rect -16 2508 83 2556
rect 1885 2508 2012 2556
rect -16 2484 2012 2508
rect 41 2010 192 2021
rect 41 1971 54 2010
rect 178 1971 192 2010
rect 41 1964 192 1971
rect 316 1966 1003 2015
rect 1094 1967 1806 2019
rect 1894 2010 2157 2020
rect 1894 1972 2031 2010
rect 2125 1972 2157 2010
rect 1894 1967 2157 1972
rect -3 1501 2025 1518
rect -3 1453 32 1501
rect 1834 1453 2025 1501
rect -3 1427 2025 1453
<< via1 >>
rect 54 1971 178 2010
rect 2031 1972 2125 2010
<< metal2 >>
rect 40 2020 2147 2022
rect 40 2010 2157 2020
rect 40 1971 54 2010
rect 178 1972 2031 2010
rect 2125 1972 2157 2010
rect 178 1971 2157 1972
rect 40 1967 2157 1971
rect 40 1962 2147 1967
use inv_module  x1
timestamp 1728978907
transform 1 0 53 0 1 1306
box -55 128 368 1254
use inv_module  x2
timestamp 1728978907
transform 1 0 844 0 1 1306
box -55 128 368 1254
use inv_module  x3
timestamp 1728978907
transform 1 0 1635 0 1 1306
box -55 128 368 1254
<< labels >>
flabel metal1 8 2513 29 2559 0 FreeSans 480 0 0 0 vdd
port 2 nsew
flabel metal1 8 1435 19 1480 0 FreeSans 480 0 0 0 gnd
port 3 nsew
flabel metal2 2141 1981 2141 1981 0 FreeSans 480 0 0 0 out
port 4 nsew
<< end >>
